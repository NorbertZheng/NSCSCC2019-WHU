module wallace_tree8_signed(a, b, z);
	/*********************
	 *	WT 8-bit Signed Multiplier
	 *input:
	 *	a[7:0]	: 8-bit 乘法器第一个操作数
	 *	b[7:0]	: 8-bit 乘法器第二个操作数
	 *output:
	 *	z[15:0]	: 16-bit 乘法器有符号结果
	 *********************/
	input [7:0] a, b;
	output [15:0] z;
	
	reg [7:0] p[7:0];
	always@(*)
		begin
		integer i, j;
		for(i = 0;i < 7;i = i + 1)
			begin
			for(j = 0;j < 7;j = j + 1)
				begin
				p[i][j] = a[i] & [j];		// AND
				end
			end
		for(i = 0;i < 7;i = i + 1)
			begin
			p[i][7] = ~(a[i] & b[7]);		// NAND
			end
		for(j = 0;j < 7;j = j + 1)
			begin
			p[7][j] = ~(a[7] & b[j]);		// NAND
			end
		p[7][7] = a[7] & b[7];
		end
	assign z[0] = p[0][0];
	
	parameter zero = 1'b0;
	parameter one = 1'b1;		// + 1000_0001_0000_0000
	wire [2:0] s1[12:01];
	wire [2:0] c1[13:02];
	add1 fa1_12_0(.a(p[7][5]), .b(p[6][6]), .ci(p[5][7]), .s(s1[12][0]), .co(c1[13][0]));
	add1 fa1_11_0(.a(p[7][4]), .b(p[6][5]), .ci(p[5][6]), .s(s1[11][0]), .co(c1[12][0]));
	add1 fa1_10_1(.a(p[7][3]), .b(p[6][4]), .ci(p[5][5]), .s(s1[10][1]), .co(c1[11][1]));
	add1 fa1_10_0(.a(p[4][6]), .b(p[3][7]), .ci(zero), .s(s1[10][0]), .co(c1[11][0]));
	add1 fa1_09_1(.a(p[7][2]), .b(p[6][3]), .ci(p[5][4]), .s(s1[09][1]), .co(c1[10][1]));
	add1 fa1_09_0(.a(p[4][5]), .b(p[3][6]), .ci(p[2][7]), .s(s1[09][0]), .co(c1[10][0]));
	add1 fa1_08_2(.a(p[7][1]), .b(p[6][2]), .ci(p[5][3]), .s(s1[08][2]), .co(c1[09][2]));
	add1 fa1_08_1(.a(p[4][4]), .b(p[3][5]), .ci(p[2][6]), .s(s1[08][1]), .co(c1[09][1]));
	add1 fa1_08_0(.a(p[1][7]), .b(one), .ci(zero), .s(s1[08][0]), .co(c1[09][0]));		// 1
	add1 fa1_07_2(.a(p[7][0]), .b(p[6][1]), .ci(p[5][2]), .s(s1[07][2]), .co(c1[08][2]));
	add1 fa1_07_1(.a(p[4][3]), .b(p[3][4]), .ci(p[2][5]), .s(s1[07][1]), .co(c1[08][1]));
	add1 fa1_07_0(.a(p[1][6]), .b(p[0][7]), .ci(zero), .s(s1[07][0]), .co(c1[08][0]));
	add1 fa1_06_1(.a(p[6][0]), .b(p[5][1]), .ci(p[4][2]), .s(s1[06][1]), .co(c1[07][1]));
	add1 fa1_06_0(.a(p[3][3]), .b(p[2][4]), .ci(p[1][5]), .s(s1[06][0]), .co(c1[07][0]));
	add1 fa1_05_1(.a(p[5][0]), .b(p[4][1]), .ci(p[3][2]), .s(s1[05][1]), .co(c1[06][1]));
	add1 fa1_05_0(.a(p[2][3]), .b(p[1][4]), .ci(p[0][5]), .s(s1[05][0]), .co(c1[06][0]));
	add1 fa1_04_1(.a(p[4][0]), .b(p[3][1]), .ci(p[2][2]), .s(s1[04][1]), .co(c1[05][1]));
	add1 fa1_04_0(.a(p[1][3]), .b(p[0][4]), .ci(zero), .s(s1[04][0]), .co(c1[05][0]));
	add1 fa1_03_0(.a(p[3][0]), .b(p[2][1]), .ci(p[1][2]), .s(s1[03][0]), .co(c1[04][0]));
	add1 fa1_02_0(.a(p[2][0]), .b(p[1][1]), .ci(p[0][2]), .s(s1[02][0]), .co(c1[03][0]));
	add1 fa1_01_0(.a(p[1][0]), .b(p[0][1]), .ci(zero), .s(s1[01][0]), .co(c1[02][0]));
	assign z[1] = s1[01][0];
	
	wire [1:0] s2[13:02];
	wire [1:0] c2[14:03];
	add1 fa2_13_0(.a(p[7][6]), .b(p[6][7]), .ci(c1[13][0]), .s(s2[13][0]), .co(c2[14][0]));
	add1 fa2_12_0(.a(s1[12][0]), .b(c1[12][0]), .ci(zero), .s(s2[12][0]), .co(c2[13][0]));
	add1 fa2_11_0(.a(s1[11][0]), .b(p[4][7]), .ci(c1[11][1]), .s(s2[11][0]), .co(c2[12][0]));
	add1 fa2_10_0(.a(s1[10][1]), .b(s1[10][0]), .ci(c1[10][1]), .s(s2[10][0]), .co(c2[11][0]));
	add1 fa2_09_1(.a(s1[09][1]), .b(s1[09][0]), .ci(c1[09][2]), .s(s2[09][1]), .co(c2[10][1]));
	add1 fa2_09_0(.a(c1[09][1]), .b(c1[09][0]), .ci(zero), .s(s2[09][0]), .co(c2[10][0]));
	add1 fa2_08_1(.a(s1[08][2]), .b(s1[08][1]), .ci(s1[08][0]), .s(s2[08][1]), .co(c2[09][1]));
	add1 fa2_08_0(.a(c1[08][2]), .b(c1[08][1]), .ci(c1[08][0]), .s(s2[08][0]), .co(c2[09][0]));
	add1 fa2_07_1(.a(s1[07][2]), .b(s1[07][1]), .ci(s1[07][0]), .s(s2[07][1]), .co(c2[08][1]));
	add1 fa2_07_0(.a(c1[07][1]), .b(c1[07][0]), .ci(zero), .s(s2[07][0]), .co(c2[08][0]));
	add1 fa2_06_1(.a(s1[06][1]), .b(s1[06][0]), .ci(p[0][6]), .s(s2[06][1]), .co(c2[07][1]));
	add1 fa2_06_0(.a(c1[06][1]), .b(c1[06][0]), .ci(zero), .s(s2[06][0]), .co(c2[07][0]));
	add1 fa2_05_0(.a(s1[05][1]), .b(s1[05][0]), .ci(c1[05][1]), .s(s2[05][0]), .co(c2[06][0]));
	add1 fa2_04_0(.a(s1[04][1]), .b(s1[04][0]), .ci(c1[04][0]), .s(s2[04][0]), .co(c2[05][0]));
	add1 fa2_03_0(.a(s1[03][0]), .b(p[0][3]), .ci(c1[03][0]), .s(s2[03][0]), .co(c2[04][0]));
	add1 fa2_02_0(.a(s1[02][0]), .b(c1[02][0]), .ci(zero), .s(s2[02][0]), .co(c2[03][0]));
	assign z[2] = s2[02][0];
	
	wire [11:03] s3;
	wire [12:04] c3;
	add1 fa3_11_0(.a(s2[11][0]), .b(c1[11][0]), .ci(c2[11][0]), .s(s3[11]), .co(c3[12]));
	add1 fa3_10_0(.a(s2[10][0]), .b(c1[10][0]), .ci(c2[10][1]), .s(s3[10]), .co(c3[11]));
	add1 fa3_09_0(.a(s2[09][1]), .b(s2[09][0]), .ci(c2[09][1]), .s(s3[09]), .co(c3[10]))
	add1 fa3_08_0(.a(s2[08][1]), .b(s2[08][0]), .ci(c2[08][1]), .s(s3[08]), .co(c3[09]));
	add1 fa3_07_0(.a(s2[07][1]), .b(s2[07][0]), .ci(c2[07][1]), .s(s3[07]), .co(c3[08]));
	add1 fa3_06_0(.a(s2[06][1]), .b(s2[06][0]), .ci(c2[06][0]), .s(s3[06]), .co(c3[07]));
	add1 fa3_05_0(.a(s2[05][0]), .b(c1[05][0]), .ci(c2[05][0]), .s(s3[05]), .co(c3[06]));
	add1 fa3_04_0(.a(s2[04][0]), .b(c2[04][0]), .ci(zero), .s(s3[04]), .co(c3[05]));
	add1 fa3_03_0(.a(s2[03][0]), .b(c2[03][0]), .ci(zero), .s(s3[03]), .co(c3[04]));
	assign z[3] = s3[03];
	
	wire [14:04] s4;
	wire [15:05] c4;
	add1 fa4_14_0(.a(p[7][7]), .b(c2[14][0]), .ci(zero), .s(s4[14]), .co(c4[15]));
	add1 fa4_13_0(.a(s2[13][0]), .b(c2[13][0]), .ci(zero), .s(s4[13]), .co(c4[14]));
	add1 fa4_12_0(.a(s2[12][0]), .b(c2[12][0]), .ci(c3[12]), .s(s4[12]), .co(c4[13]));
	add1 fa4_11_0(.a(s3[11]), .b(c3[11]), .ci(zero), .s(s4[11]), .co(c4[12]));
	add1 fa4_10_0(.a(s3[10]), .b(c2[10][0]), .ci(c3[10]), .s(s4[10]), .co(c4[11]));
	add1 fa4_09_0(.a(s3[09]), .b(c2[09][0]), .ci(c3[09]), .s(s4[09]), .co(c4[10]));
	add1 fa4_08_0(.a(s3[08]), .b(c2[08][0]), .ci(c3[08]), .s(s4[08]), .co(c4[09]));
	add1 fa4_07_0(.a(s3[07]), .b(c2[07][0]), .ci(c3[07]), .s(s4[07]), .co(c4[08]));
	add1 fa4_06_0(.a(s3[06]), .b(c3[06]), .ci(zero), .s(s4[06]), .co(c4[07]));
	add1 fa4_05_0(.a(s3[05]), .b(c3[05]), .ci(zero), .s(s4[05]), .co(c4[06]));
	add1 fa4_04_0(.a(s3[04]), .b(c3[04]), .ci(zero), .s(s4[04]), .co(c4[05]));
	assign z[4] = s4[04];
	
	assign z[15:5] = {one, s4[14:05]} + c4[15:05];		// 1
endmodule